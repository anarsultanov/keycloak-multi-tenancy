dev.sultanov.keycloak.multitenancy.model.TenantSpi